module arrow(input logic [9:0] addr,
				output logic [0:99]data);
					
parameter stand_width = 100;
parameter stand_lenth = 100;


parameter [0:stand_lenth-1][0:stand_width-1] ROM = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000000011111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000000011111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
};
assign data = ROM[addr][0:99];
endmodule


					