module kick(input logic [9:0] addr,
				input logic frame_clk,  kick,
				output logic kick_1, kick_valid,
					 output logic [0:99]data);
		  
enum logic [2:0] {stand, kick1, kick2, Wait}state, next_state;		
logic [4:0] counter, counter1; 
parameter stand_width = 100;
parameter stand_lenth = 100;


parameter [0:stand_lenth-1][0:stand_width-1] ROM = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111000000011000001000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000010000001100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000110000001100000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000001110000001110000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000001110000011111000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000011110000011111000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000111110000011111100000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000111110000011111110000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111110000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111100000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111100000001111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111110000000111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111000000000001111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111000000000000111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111110000000000111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111100000011111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111001111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000001111000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000111100000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
};

parameter [0:stand_lenth-1][0:stand_width-1] ROM1 = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000011000001000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111000000010000001100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111000000110000001100000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000001110000001110000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000001110000011111000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000011110000011111000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000111110000011111100000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000111110000011111110000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111110000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111100000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111100000001111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111110000000111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111000000000001111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111000000000000111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111110000000000111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111100000011111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000111111100000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111001111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001100000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001110000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111100000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111100000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111110000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111000000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111000000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111100000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111110000000111111111000111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111000000011111110000011111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111100000011111100000011111111111111111,
100'b1111111111111111111111111111111111111111111100000111111111111111110000001111000000011111111111111111,
100'b1111111111111111111111111111111111111111111000000111111111111111110000000110000000011111111111111111,
100'b1111111111111111111111111111111111111111111000000111111111111111111000000000000000111111111111111111,
100'b1111111111111111111111111111111111111111111000001111111111111111111100000000000001111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111100000000000111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111110000000001111111111111111111111,
100'b1111111111111111111111111111111111111111110000011111111111111111111110000000011111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111000000111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
};

parameter [0:stand_lenth-1][0:stand_width-1] ROM2 = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111111100001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111111000000111111111111111000001111111111111111,
100'b1111111111111111111111111111111111111111000000011111111111000000111111111111110000000011111111111111,
100'b1111111111111111111111111111111111111110000000001111111110000001111111111111110000000001111111111111,
100'b1111111111111111111111111111111111111100000000000111111100000001111111111111110000000000111111111111,
100'b1111111111111111111111111111111111111000000000000011111100000011111111111111111100000000111111111111,
100'b1111111111111111111111111111111111111000000000000011111100000111111111111111111110000000011111111111,
100'b1111111111111111111111111111111111110000000000000001111000000111111111111111111100000000011111111111,
100'b1111111111111111111111111111111111110000000000000000111000001111111111111111111000000000111111111111,
100'b1111111111111111111111111111111111100000000000000000111000001111111111111111110000000001111111111111,
100'b1111111111111111111111111111111111100000000000000000110000011111111111111111000000000011111111111111,
100'b1111111111111111111111111111111111100000000000000000010000011111111111111110000000001111111111111111,
100'b1111111111111111111111111111111111000000110000010000000000011111111111111100000000011111111111111111,
100'b1111111111111111111111111111111111000000110000011000000000011111111111111000000001111111111111111111,
100'b1111111111111111111111111111111110000001110000011000000000111111111111100000000011111111111111111111,
100'b1111111111111111111111111111111110000001110000011100000001111111111111000000000111111111111111111111,
100'b1111111111111111111111111111111100000011110000011100000001111111111100000000011111111111111111111111,
100'b1111111111111111111111111111111100000011110000001100000011111111111000000000111111111111111111111111,
100'b1111111111111111111111111111111100000111111000001110000111111111110000000011111111111111111111111111,
100'b1111111111111111111111111111111000000111111000001111111111111111000000000111111111111111111111111111,
100'b1111111111111111111111111111111000000111111000001111111111111110000000001111111111111111111111111111,
100'b1111111111111111111111111111110000001111111000000111111111111000000000111111111111111111111111111111,
100'b1111111111111111111111111111110000001111111000000111111111110000000001111111111111111111111111111111,
100'b1111111111111111111111111111110000001111111100000111111111000000000011111111111111111111111111111111,
100'b1111111111111111111111111111110000001111111100000011111110000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111000000111111100000001111000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111000000111111100000000100000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000111111110000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000111111110000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000011111110000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111100000011111111000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000111111111000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111001111111111000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
};


always_ff @(posedge frame_clk) begin
	state <= next_state;
	if(counter == 5'd10) 
		counter <= 5'b0;
	else 
		counter <= counter + 1'b1;
		
	if(counter1 == 5'd29) 
		counter1 <= 5'b0;
	else 
		counter1 <= counter1 + 1'b1;
	end
	
always_comb 
	begin
	next_state = state;
		case(state) 
		stand:
			if(counter == 5'd9 && kick)
			next_state = kick1;
			else 
			next_state = stand;
		kick1:
			if(counter == 5'd9)
			next_state = kick2;
			else
			next_state = kick1;
		kick2:
			if(counter == 5'd9)
			next_state = Wait;
			else
			next_state = kick2;
		Wait:
			if(counter1 == 5'd28)
			next_state = stand;
			else 
			next_state = Wait;
			
		endcase
	end

always_comb 
	begin
	data = data;
	kick_1 = kick_1;
	kick_valid = kick_valid;
		case(state) 
		stand: 	begin
			data = ROM[addr][0:99];
			kick_1 = 1'b0;
			kick_valid = 1'b0;
				end

		kick1:	begin
			data = ROM1[addr][0:99];
			kick_1 = 1'b1;
			kick_valid = 1'b0;
				end
				
		kick2:	begin
			data = ROM2[addr][0:99];
			kick_1 = 1'b1;
			kick_valid = 1'b1;
				end
		Wait: begin
			data = ROM[addr][0:99];
			kick_1 = 1'b0;
			kick_valid = 1'b0;
				end
			
					
		endcase
	end

	
	

endmodule 