module jump(input logic [9:0] addr,
					 input logic jump, frame_clk,
					 output logic jump_1, jump_valid,
					 output logic [0:99]data);
		  
enum logic [2:0] {stand, jump1, jump2, jump3, jump4, Wait} state, next_state;		
logic [4:0] counter, counter1; 
parameter stand_width = 100;
parameter stand_lenth = 100;


parameter [0:stand_lenth-1][0:stand_width-1] ROM = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111000000011000001000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000010000001100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000110000001100000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000001110000001110000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000001110000011111000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000011110000011111000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000111110000011111100000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000111110000011111110000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111110000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111100000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111100000001111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111110000000100001111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111000000000001111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111000000000000111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111110000000000111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111100000011111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111001111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000001111000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000111100000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
};

parameter [0:stand_lenth-1][0:stand_width-1] ROM1 = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000001111001111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000001110000111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000001110000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000000001100000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000000001100000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000000001100000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001000001100000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000010000001100000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001100000001100000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001000000011100000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000011000000011000000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000010000000000000000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000000000000000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111100011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111110000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111100000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011110000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011110000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111100000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111000000010000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111000000110000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000010000001110000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000001110000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000001111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000011111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000111111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000001111111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000001111111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111000000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111000000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111100000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111110000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111111110111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111};

parameter [0:stand_lenth-1][0:stand_width-1] ROM2 = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000010000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000010000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000000000000111111111111000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000000000000111111111100000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000000000000111111110000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000000000000011110000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000000000000011000000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000000000000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000100000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000100000000001110000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111001110000000001100000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111110000000000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111};

parameter [0:stand_lenth-1][0:stand_width-1] ROM3 = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000100000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111100000000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000111111000000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000111111100000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000011111110000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000100000011111110000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001100000011111110000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000001100000011111100000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011100000011111100000011111111111111111111111111111111,
100'b1111111111111111111111111111111000000000000000111100000011111100000111111111111111111111111111111111,
100'b1111111111111111111111111111110000000000000000111100000011111100000111111111111111111111111111111111,
100'b1111111111111111111111111111110000000000000001111100000011111100000111111111111111111111111111111111,
100'b1111111111111111111111111111110000000000000011111110000011111100001111111111111111111111111111111111,
100'b1111111111111111111111111111111000000000000111111110000011111100001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000001111111001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000001110000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000001111000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000011111000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000110000001111000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000000111110111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111};

parameter [0:stand_lenth-1][0:stand_width-1] ROM4 = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000111110011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000011100001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000001000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111001111111111000000000000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000111111111000000000000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111111000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111110000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111110000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111000001111100000000000010000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111000001111000000000000011000000001111111111111111100011111111111111,
100'b1111111111111111111111111111111111000000111000000100000011100000001111111111111111000000001111111111,
100'b1111111111111111111111111111111111000000110000001100000011110000000111111111111111000000000011111111,
100'b1111111111111111111111111111111111100000000000001100000011110000000111111111111111000000000001111111,
100'b1111111111111111111111111111111111100000000000011100000011111000000111111111111111000000000001111111,
100'b1111111111111111111111111111111111110000000000111100000011111000000111111111111110000000000001111111,
100'b1111111111111111111111111111111111110000000000111100000011111100001111111111111000000000000011111111,
100'b1111111111111111111111111111111111111000000001111100000011111111111111111111000000000000000111111111,
100'b1111111111111111111111111111111111111100000111111110000011111111111111111000000000000001111111111111,
100'b1111111111111111111111111111111111111110001111111110000011111111111111100000000000000111111111111111,
100'b1111111111111111111111111111111111111111111111111110000011111111111100000000000000011111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111110000000000000001111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111000000000000001111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111000000000000001111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001000000000000000111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111101100000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111};

always_ff @(posedge frame_clk) begin
	state <= next_state;
	if(counter == 5'd10) 
		counter <= 5'b0;
	else 
		counter <= counter + 1'b1;
	
	if(counter1 == 5'd29) 
		counter1 <= 5'b0;
	else 
		counter1 <= counter1 + 1'b1;
	end
	
always_comb 
	begin
	next_state = state;
		case(state) 
		stand:
			if(counter == 5'd9 && jump)
			next_state = jump1;
			else 
			next_state = stand;
		jump1:
			if(counter == 5'd9)
			next_state = jump2;
			else
			next_state = jump1;
		jump2:
			if(counter == 5'd9)
			next_state = jump3;
			else
			next_state = jump2;
		jump3:
			if(counter == 5'd9)
			next_state = jump4;
			else
			next_state = jump3;
		jump4:
			if(counter == 5'd9)
			next_state = Wait;
			else
			next_state = jump4;
		Wait:
			if(counter1 == 5'd28)
			next_state = stand;
			else 
			next_state = Wait;
		endcase
	end

always_comb 
	begin
	data = data;
	jump_1 = jump_1;
	jump_valid = jump_valid;
	
		case(state) 
		stand: begin
			data = ROM[addr][0:99];
			jump_1 = 1'b0;
			jump_valid = 1'b0;
				end
		jump1:	begin
			data = ROM1[addr][0:99];
				jump_1 = 1'b1;
				jump_valid = 1'b0;
				end
		jump2:	begin
			data = ROM2[addr][0:99];
				jump_1 = 1'b1;
				jump_valid = 1'b0;
				end
		jump3:	begin
			data = ROM3[addr][0:99];
				jump_1 = 1'b1;
				jump_valid = 1'b0;
				end
		jump4:	begin
			data = ROM4[addr][0:99];
				jump_1 = 1'b1;
				jump_valid = 1'b1;
				end
		Wait: begin
			data = ROM[addr][0:99];
			jump_1 = 1'b0;
			jump_valid = 1'b0;
				end
		endcase
	end

	
	

endmodule 