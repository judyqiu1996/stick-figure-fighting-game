module back(input logic [9:0] addr,
					input logic frame_clk, back, Clk,
					output logic back_1, 
					 output logic [0:99]data);
		  
enum logic [2:0] {stand, back1, back2}state, next_state;		
logic [4:0] counter;
logic [5:0] counter1; 
parameter stand_width = 100;
parameter stand_lenth = 100;


parameter [0:stand_lenth-1][0:stand_width-1] ROM = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111000000011000001000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000010000001100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000110000001100000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000001110000001110000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111100000001110000011111000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000011110000011111000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000111110000011111100000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000111110000011111110000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111110000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111100000011111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111100000001111111111111111111111111111111111,
100'b1111111111111111111111111111111110000001111100000011111111110000000111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111000000000001111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111000000000000111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000011111111111110000000000111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111100000011111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000011111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111001111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000001111000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000111100000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
};

parameter [0:stand_lenth-1][0:stand_width-1] ROM1 = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000001111111111000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000001111111110000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000111111110000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000000111111100000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111100000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111100000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000000111000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000000000000111000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000110000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000000000000100000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000110000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000011111000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000011111100000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000000011111110000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000001111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000001000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011100000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111110000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111110000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000111111111000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000001111000000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000000000111000000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000000111100000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000000001111111111110011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,

};

parameter [0:stand_lenth-1][0:stand_width-1] ROM2 = {
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111000011111110000001111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111000001110000000000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111000001100000000000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111100111111100000000000000000000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111000001111110000000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111110000000111110000000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111000000011110000000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111000000001110000000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111100000001110000000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111110000000110000000000000000000000001111111111111111111111111111111111111111111111,
100'b1111111111111111111111000000011000000000000000000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111100000001000000000000000000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111110000001000000000000000000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111110000000100000000000000000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111000000010000000000000000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111100000011000000000000000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111100000001100000000000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111110000000100000000000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111000000010000000001111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111110000000100000000011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000110000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111000000011000000000011111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111100000011110000000001111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000001111000000000111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111110000001111110000000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111000000111111000000011111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111000000111111100000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111110000001111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111100000011111111000000111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111110000001111111000000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111110000001111111100000011111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111000001111111110000001111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111000000111111110000001111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111000000111111111000000111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000111111111000000111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000011111111100000011111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111100000011111111100000011111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000011111111110000000000111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000011111111110000000000111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000001111111111000000000111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000001111111111000000000111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111110000001111111111100000001111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111000001111111111110001111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111

};


always_ff @(posedge frame_clk) begin
	state <= next_state;
	if(counter == 5'd10) 
		counter <= 5'b0;
	else 
		counter <= counter + 1'b1;
		
	if(counter1 == 6'd40) 
		counter1 <= 6'b0;
	else 
		counter1 <= counter1 + 1'b1;
	end
	
always_comb 
	begin
	next_state = state;
		case(state) 
		stand:
			if(back)
			next_state = back1;
			else 
			next_state = stand;
		back1:
			if(counter == 5'd9)
			next_state = back2;
			else
			next_state = back1;
		back2:
			if(counter1 == 6'd39 && ~back)
			next_state = stand;
			else
			next_state = back2;

		endcase
	end

always_comb 
	begin
			data = 0;
			back_1 = 0;

		case(state) 
		
		stand: begin
			data = ROM[addr][0:99];
			back_1 = 1'b0;
				end

		back1:	begin
			data = ROM1[addr][0:99];
			back_1 =1'b1;
			end

		back2:	begin
			data = ROM2[addr][0:99];
			back_1 =1'b1;
					end

		endcase
	end

	
	

endmodule 