module collision(input logic near0, stand_right, stand_left, attck, 
					  input logic [9:0]positionX, positionY, positionX1, positionY1,
					  output logic valid);
					  
	if (near0 )
					  
	